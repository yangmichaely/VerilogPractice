module queue(
    input wire [31:0] in,
    input signal,
    output wire [31:0] out,
    output queue_full,
    output queue_empty
);

