module hw4_tb();

int test_num;
reg 